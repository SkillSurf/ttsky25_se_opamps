magic
tech sky130A
magscale 1 2
timestamp 1591351771
<< checkpaint >>
rect -3732 -3932 34474 49084
<< metal1 >>
rect 200 41534 600 41568
rect 200 41533 325 41534
rect 200 41481 238 41533
rect 290 41482 325 41533
rect 377 41482 422 41534
rect 474 41482 502 41534
rect 554 41482 600 41534
rect 290 41481 600 41482
rect 200 41454 600 41481
rect 200 41453 325 41454
rect 200 41401 238 41453
rect 290 41402 325 41453
rect 377 41402 422 41454
rect 474 41402 502 41454
rect 554 41402 600 41454
rect 290 41401 600 41402
rect 200 41368 600 41401
rect 20734 41541 20914 41556
rect 20734 41489 20758 41541
rect 20810 41489 20838 41541
rect 20890 41489 20914 41541
rect 20734 41461 20914 41489
rect 20734 41409 20758 41461
rect 20810 41409 20838 41461
rect 20890 41409 20914 41461
rect 20734 41392 20914 41409
rect 2756 24314 2936 24329
rect 2756 24262 2780 24314
rect 2832 24262 2860 24314
rect 2912 24262 2936 24314
rect 2756 24234 2936 24262
rect 2756 24182 2780 24234
rect 2832 24182 2860 24234
rect 2912 24182 2936 24234
rect 2756 24165 2936 24182
rect 2162 23659 2342 23674
rect 2162 23607 2186 23659
rect 2238 23607 2266 23659
rect 2318 23607 2342 23659
rect 2162 23579 2342 23607
rect 2162 23527 2186 23579
rect 2238 23527 2266 23579
rect 2318 23527 2342 23579
rect 2162 23510 2342 23527
rect 2162 18252 2262 23510
rect 2756 18457 2856 24165
rect 2162 18152 2755 18252
rect 5557 10738 6143 10740
rect 5557 10686 5851 10738
rect 5903 10686 5915 10738
rect 5967 10686 6007 10738
rect 6059 10686 6071 10738
rect 6123 10686 6143 10738
rect 5557 10684 6143 10686
rect 5557 7174 5616 10684
<< via1 >>
rect 238 41481 290 41533
rect 325 41482 377 41534
rect 422 41482 474 41534
rect 502 41482 554 41534
rect 238 41401 290 41453
rect 325 41402 377 41454
rect 422 41402 474 41454
rect 502 41402 554 41454
rect 20758 41489 20810 41541
rect 20838 41489 20890 41541
rect 20758 41409 20810 41461
rect 20838 41409 20890 41461
rect 2780 24262 2832 24314
rect 2860 24262 2912 24314
rect 2780 24182 2832 24234
rect 2860 24182 2912 24234
rect 2186 23607 2238 23659
rect 2266 23607 2318 23659
rect 2186 23527 2238 23579
rect 2266 23527 2318 23579
rect 11818 17669 11870 17721
rect 11898 17669 11950 17721
rect 11818 17589 11870 17641
rect 11898 17589 11950 17641
rect 5851 10686 5903 10738
rect 5915 10686 5967 10738
rect 6007 10686 6059 10738
rect 6071 10686 6123 10738
rect 1897 10494 1949 10546
rect 1897 10430 1949 10482
rect 1897 7174 1949 7226
rect 1897 7110 1949 7162
<< metal2 >>
rect 200 41536 600 41568
rect 200 41535 323 41536
rect 200 41479 236 41535
rect 292 41480 323 41535
rect 379 41480 420 41536
rect 292 41479 420 41480
rect 200 41456 420 41479
rect 200 41455 323 41456
rect 200 41399 236 41455
rect 292 41400 323 41455
rect 379 41400 420 41456
rect 556 41400 600 41536
rect 292 41399 600 41400
rect 200 41368 600 41399
rect 20734 41543 20914 41556
rect 20734 41407 20756 41543
rect 20892 41407 20914 41543
rect 20734 41392 20914 41407
rect 3026 39988 3114 41347
rect 2735 39900 3114 39988
rect 2735 25055 2823 39900
rect 3036 25959 3124 38901
rect 26451 37617 26618 37630
rect 26451 37526 26468 37617
rect 19458 37481 26468 37526
rect 26604 37481 26618 37617
rect 19458 37466 26618 37481
rect 19549 26606 19637 35910
rect 30362 26634 30542 26647
rect 30362 26606 30384 26634
rect 19549 26518 30384 26606
rect 30362 26498 30384 26518
rect 30520 26498 30542 26634
rect 30362 26483 30542 26498
rect 26498 25984 26678 25997
rect 26498 25959 26520 25984
rect 3036 25871 26520 25959
rect 26498 25848 26520 25871
rect 26656 25848 26678 25984
rect 26498 25833 26678 25848
rect 22634 25080 22814 25093
rect 22634 25055 22656 25080
rect 2735 24967 22656 25055
rect 22634 24944 22656 24967
rect 22792 24944 22814 25080
rect 22634 24929 22814 24944
rect 27003 24420 27170 24433
rect 27003 24329 27020 24420
rect 2756 24314 27020 24329
rect 2756 24262 2780 24314
rect 2832 24262 2860 24314
rect 2912 24284 27020 24314
rect 27156 24284 27170 24420
rect 2912 24269 27170 24284
rect 2912 24262 2936 24269
rect 2756 24234 2936 24262
rect 2756 24182 2780 24234
rect 2832 24182 2860 24234
rect 2912 24182 2936 24234
rect 2756 24165 2936 24182
rect 30362 23697 30542 23710
rect 30362 23674 30384 23697
rect 2162 23659 30384 23674
rect 2162 23607 2186 23659
rect 2238 23607 2266 23659
rect 2318 23607 30384 23659
rect 2162 23582 30384 23607
rect 2162 23579 2342 23582
rect 2162 23527 2186 23579
rect 2238 23527 2266 23579
rect 2318 23527 2342 23579
rect 30362 23561 30384 23582
rect 30520 23561 30542 23697
rect 30362 23546 30542 23561
rect 2162 23510 2342 23527
rect 200 22605 2724 22637
rect 200 22604 323 22605
rect 200 22548 236 22604
rect 292 22549 323 22604
rect 379 22549 420 22605
rect 292 22548 420 22549
rect 200 22525 420 22548
rect 200 22524 323 22525
rect 200 22468 236 22524
rect 292 22469 323 22524
rect 379 22469 420 22525
rect 556 22469 2724 22605
rect 292 22468 2724 22469
rect 200 22437 2724 22468
rect 1252 19554 2460 19618
rect 1252 14430 1352 19554
rect 1426 19383 2460 19447
rect 1426 15117 1526 19383
rect 11794 17723 11974 17736
rect 11794 17587 11816 17723
rect 11952 17587 11974 17723
rect 11794 17572 11974 17587
rect 1601 17195 1960 17223
rect 1601 17194 1705 17195
rect 1601 17138 1618 17194
rect 1674 17139 1705 17194
rect 1761 17139 1802 17195
rect 1674 17138 1802 17139
rect 1601 17115 1802 17138
rect 1601 17114 1705 17115
rect 1601 17058 1618 17114
rect 1674 17059 1705 17114
rect 1761 17059 1802 17115
rect 1938 17059 1960 17195
rect 1674 17058 1960 17059
rect 1601 17031 1960 17058
rect 22634 15138 22814 15151
rect 22634 15117 22656 15138
rect 1426 15017 22656 15117
rect 22634 15002 22656 15017
rect 22792 15002 22814 15138
rect 22634 14987 22814 15002
rect 26498 14451 26678 14464
rect 26498 14430 26520 14451
rect 1252 14330 26520 14430
rect 26498 14315 26520 14330
rect 26656 14315 26678 14451
rect 26498 14300 26678 14315
rect 200 13323 6256 13378
rect 200 13322 323 13323
rect 200 13266 236 13322
rect 292 13267 323 13322
rect 379 13267 420 13323
rect 292 13266 420 13267
rect 200 13243 420 13266
rect 200 13242 323 13243
rect 200 13186 236 13242
rect 292 13187 323 13242
rect 379 13187 420 13243
rect 556 13187 6256 13323
rect 292 13186 6256 13187
rect 200 13130 6256 13186
rect 18770 13000 18950 13013
rect 18770 12959 18792 13000
rect 8466 12903 18792 12959
rect 18770 12864 18792 12903
rect 18928 12864 18950 13000
rect 18770 12849 18950 12864
rect 22634 10784 22814 10797
rect 22634 10740 22656 10784
rect 5831 10738 22656 10740
rect 5831 10686 5851 10738
rect 5903 10686 5915 10738
rect 5967 10686 6007 10738
rect 6059 10686 6071 10738
rect 6123 10686 22656 10738
rect 5831 10684 22656 10686
rect 22634 10648 22656 10684
rect 22792 10648 22814 10784
rect 22634 10633 22814 10648
rect 1895 10546 1951 10566
rect 1895 10494 1897 10546
rect 1949 10494 1951 10546
rect 1895 10482 1951 10494
rect 1895 10430 1897 10482
rect 1949 10430 1951 10482
rect 1895 7226 1951 10430
rect 1895 7174 1897 7226
rect 1949 7174 1951 7226
rect 1895 7162 1951 7174
rect 1895 7110 1897 7162
rect 1949 7110 1951 7162
rect 1895 5737 1951 7110
rect 1329 5651 1951 5737
rect 1329 1878 1428 5651
rect 5106 4685 5274 4711
rect 5106 4666 5119 4685
rect 4972 4549 5119 4666
rect 5255 4549 5274 4685
rect 4972 4519 5274 4549
rect 1460 2135 1554 4458
rect 27556 2424 27723 2437
rect 27556 2333 27573 2424
rect 5494 2288 27573 2333
rect 27709 2288 27723 2424
rect 5494 2273 27723 2288
rect 30362 2158 30542 2171
rect 30362 2135 30384 2158
rect 1460 2043 30384 2135
rect 30362 2022 30384 2043
rect 30520 2022 30542 2158
rect 30362 2007 30542 2022
rect 26498 1901 26678 1914
rect 26498 1878 26520 1901
rect 1329 1784 26520 1878
rect 26498 1765 26520 1784
rect 26656 1765 26678 1901
rect 26498 1750 26678 1765
<< via2 >>
rect 236 41533 292 41535
rect 236 41481 238 41533
rect 238 41481 290 41533
rect 290 41481 292 41533
rect 236 41479 292 41481
rect 323 41534 379 41536
rect 323 41482 325 41534
rect 325 41482 377 41534
rect 377 41482 379 41534
rect 323 41480 379 41482
rect 420 41534 556 41536
rect 420 41482 422 41534
rect 422 41482 474 41534
rect 474 41482 502 41534
rect 502 41482 554 41534
rect 554 41482 556 41534
rect 236 41453 292 41455
rect 236 41401 238 41453
rect 238 41401 290 41453
rect 290 41401 292 41453
rect 236 41399 292 41401
rect 323 41454 379 41456
rect 323 41402 325 41454
rect 325 41402 377 41454
rect 377 41402 379 41454
rect 323 41400 379 41402
rect 420 41454 556 41482
rect 420 41402 422 41454
rect 422 41402 474 41454
rect 474 41402 502 41454
rect 502 41402 554 41454
rect 554 41402 556 41454
rect 420 41400 556 41402
rect 20756 41541 20892 41543
rect 20756 41489 20758 41541
rect 20758 41489 20810 41541
rect 20810 41489 20838 41541
rect 20838 41489 20890 41541
rect 20890 41489 20892 41541
rect 20756 41461 20892 41489
rect 20756 41409 20758 41461
rect 20758 41409 20810 41461
rect 20810 41409 20838 41461
rect 20838 41409 20890 41461
rect 20890 41409 20892 41461
rect 20756 41407 20892 41409
rect 26468 37481 26604 37617
rect 30384 26498 30520 26634
rect 26520 25848 26656 25984
rect 22656 24944 22792 25080
rect 27020 24284 27156 24420
rect 30384 23561 30520 23697
rect 236 22548 292 22604
rect 323 22549 379 22605
rect 236 22468 292 22524
rect 323 22469 379 22525
rect 420 22469 556 22605
rect 11816 17721 11952 17723
rect 11816 17669 11818 17721
rect 11818 17669 11870 17721
rect 11870 17669 11898 17721
rect 11898 17669 11950 17721
rect 11950 17669 11952 17721
rect 11816 17641 11952 17669
rect 11816 17589 11818 17641
rect 11818 17589 11870 17641
rect 11870 17589 11898 17641
rect 11898 17589 11950 17641
rect 11950 17589 11952 17641
rect 11816 17587 11952 17589
rect 1618 17138 1674 17194
rect 1705 17139 1761 17195
rect 1618 17058 1674 17114
rect 1705 17059 1761 17115
rect 1802 17059 1938 17195
rect 22656 15002 22792 15138
rect 26520 14315 26656 14451
rect 236 13266 292 13322
rect 323 13267 379 13323
rect 236 13186 292 13242
rect 323 13187 379 13243
rect 420 13187 556 13323
rect 18792 12864 18928 13000
rect 22656 10648 22792 10784
rect 5119 4549 5255 4685
rect 27573 2288 27709 2424
rect 30384 2022 30520 2158
rect 26520 1765 26656 1901
<< metal3 >>
rect 219 41540 578 41564
rect 219 41539 319 41540
rect 219 41475 232 41539
rect 296 41476 319 41539
rect 383 41476 416 41540
rect 296 41475 416 41476
rect 219 41460 416 41475
rect 219 41459 319 41460
rect 219 41395 232 41459
rect 296 41396 319 41459
rect 383 41396 416 41460
rect 560 41396 578 41540
rect 296 41395 578 41396
rect 219 41372 578 41395
rect 20734 41547 20914 41556
rect 20734 41403 20752 41547
rect 20896 41403 20914 41547
rect 20734 41392 20914 41403
rect 26451 37621 26618 37630
rect 26451 37477 26464 37621
rect 26608 37477 26618 37621
rect 26451 37466 26618 37477
rect 2106 33765 2465 33789
rect 2106 33764 2206 33765
rect 2106 33700 2119 33764
rect 2183 33701 2206 33764
rect 2270 33701 2303 33765
rect 2183 33700 2303 33701
rect 2106 33685 2303 33700
rect 2106 33684 2206 33685
rect 2106 33620 2119 33684
rect 2183 33621 2206 33684
rect 2270 33621 2303 33685
rect 2447 33621 2465 33765
rect 2183 33620 2465 33621
rect 2106 33597 2465 33620
rect 30362 26638 30542 26647
rect 30362 26494 30380 26638
rect 30524 26494 30542 26638
rect 30362 26483 30542 26494
rect 26498 25988 26678 25997
rect 26498 25844 26516 25988
rect 26660 25844 26678 25988
rect 26498 25833 26678 25844
rect 22634 25084 22814 25093
rect 22634 24940 22652 25084
rect 22796 24940 22814 25084
rect 22634 24929 22814 24940
rect 27003 24424 27170 24433
rect 27003 24280 27016 24424
rect 27160 24280 27170 24424
rect 27003 24269 27170 24280
rect 30362 23701 30542 23710
rect 30362 23557 30380 23701
rect 30524 23557 30542 23701
rect 30362 23546 30542 23557
rect 219 22609 578 22633
rect 219 22608 319 22609
rect 219 22544 232 22608
rect 296 22545 319 22608
rect 383 22545 416 22609
rect 296 22544 416 22545
rect 219 22529 416 22544
rect 219 22528 319 22529
rect 219 22464 232 22528
rect 296 22465 319 22528
rect 383 22465 416 22529
rect 560 22465 578 22609
rect 296 22464 578 22465
rect 219 22441 578 22464
rect 11794 17727 11974 17736
rect 11794 17583 11812 17727
rect 11956 17583 11974 17727
rect 11794 17572 11974 17583
rect 1601 17199 1960 17223
rect 1601 17198 1701 17199
rect 1601 17134 1614 17198
rect 1678 17135 1701 17198
rect 1765 17135 1798 17199
rect 1678 17134 1798 17135
rect 1601 17119 1798 17134
rect 1601 17118 1701 17119
rect 1601 17054 1614 17118
rect 1678 17055 1701 17118
rect 1765 17055 1798 17119
rect 1942 17055 1960 17199
rect 1678 17054 1960 17055
rect 1601 17031 1960 17054
rect 22634 15142 22814 15151
rect 22634 14998 22652 15142
rect 22796 14998 22814 15142
rect 22634 14987 22814 14998
rect 26498 14455 26678 14464
rect 26498 14311 26516 14455
rect 26660 14311 26678 14455
rect 26498 14300 26678 14311
rect 219 13327 578 13351
rect 219 13326 319 13327
rect 219 13262 232 13326
rect 296 13263 319 13326
rect 383 13263 416 13327
rect 296 13262 416 13263
rect 219 13247 416 13262
rect 219 13246 319 13247
rect 219 13182 232 13246
rect 296 13183 319 13246
rect 383 13183 416 13247
rect 560 13183 578 13327
rect 296 13182 578 13183
rect 219 13159 578 13182
rect 18770 13004 18950 13013
rect 18770 12860 18788 13004
rect 18932 12860 18950 13004
rect 18770 12849 18950 12860
rect 22634 10788 22814 10797
rect 22634 10644 22652 10788
rect 22796 10644 22814 10788
rect 22634 10633 22814 10644
rect 4935 4687 5274 4711
rect 4935 4686 5035 4687
rect 4935 4622 4948 4686
rect 5012 4623 5035 4686
rect 5099 4685 5274 4687
rect 5099 4623 5119 4685
rect 5012 4622 5119 4623
rect 4935 4607 5119 4622
rect 4935 4606 5035 4607
rect 4935 4542 4948 4606
rect 5012 4543 5035 4606
rect 5099 4549 5119 4607
rect 5255 4549 5274 4685
rect 5099 4543 5274 4549
rect 5012 4542 5274 4543
rect 4935 4519 5274 4542
rect 27556 2428 27723 2437
rect 27556 2284 27569 2428
rect 27713 2284 27723 2428
rect 27556 2273 27723 2284
rect 30362 2162 30542 2171
rect 30362 2018 30380 2162
rect 30524 2018 30542 2162
rect 30362 2007 30542 2018
rect 26498 1905 26678 1914
rect 26498 1761 26516 1905
rect 26660 1761 26678 1905
rect 26498 1750 26678 1761
<< via3 >>
rect 232 41535 296 41539
rect 232 41479 236 41535
rect 236 41479 292 41535
rect 292 41479 296 41535
rect 232 41475 296 41479
rect 319 41536 383 41540
rect 319 41480 323 41536
rect 323 41480 379 41536
rect 379 41480 383 41536
rect 319 41476 383 41480
rect 416 41536 560 41540
rect 232 41455 296 41459
rect 232 41399 236 41455
rect 236 41399 292 41455
rect 292 41399 296 41455
rect 232 41395 296 41399
rect 319 41456 383 41460
rect 319 41400 323 41456
rect 323 41400 379 41456
rect 379 41400 383 41456
rect 319 41396 383 41400
rect 416 41400 420 41536
rect 420 41400 556 41536
rect 556 41400 560 41536
rect 416 41396 560 41400
rect 20752 41543 20896 41547
rect 20752 41407 20756 41543
rect 20756 41407 20892 41543
rect 20892 41407 20896 41543
rect 20752 41403 20896 41407
rect 26464 37617 26608 37621
rect 26464 37481 26468 37617
rect 26468 37481 26604 37617
rect 26604 37481 26608 37617
rect 26464 37477 26608 37481
rect 2119 33700 2183 33764
rect 2206 33701 2270 33765
rect 2119 33620 2183 33684
rect 2206 33621 2270 33685
rect 2303 33621 2447 33765
rect 30380 26634 30524 26638
rect 30380 26498 30384 26634
rect 30384 26498 30520 26634
rect 30520 26498 30524 26634
rect 30380 26494 30524 26498
rect 26516 25984 26660 25988
rect 26516 25848 26520 25984
rect 26520 25848 26656 25984
rect 26656 25848 26660 25984
rect 26516 25844 26660 25848
rect 22652 25080 22796 25084
rect 22652 24944 22656 25080
rect 22656 24944 22792 25080
rect 22792 24944 22796 25080
rect 22652 24940 22796 24944
rect 27016 24420 27160 24424
rect 27016 24284 27020 24420
rect 27020 24284 27156 24420
rect 27156 24284 27160 24420
rect 27016 24280 27160 24284
rect 30380 23697 30524 23701
rect 30380 23561 30384 23697
rect 30384 23561 30520 23697
rect 30520 23561 30524 23697
rect 30380 23557 30524 23561
rect 232 22604 296 22608
rect 232 22548 236 22604
rect 236 22548 292 22604
rect 292 22548 296 22604
rect 232 22544 296 22548
rect 319 22605 383 22609
rect 319 22549 323 22605
rect 323 22549 379 22605
rect 379 22549 383 22605
rect 319 22545 383 22549
rect 416 22605 560 22609
rect 232 22524 296 22528
rect 232 22468 236 22524
rect 236 22468 292 22524
rect 292 22468 296 22524
rect 232 22464 296 22468
rect 319 22525 383 22529
rect 319 22469 323 22525
rect 323 22469 379 22525
rect 379 22469 383 22525
rect 319 22465 383 22469
rect 416 22469 420 22605
rect 420 22469 556 22605
rect 556 22469 560 22605
rect 416 22465 560 22469
rect 11812 17723 11956 17727
rect 11812 17587 11816 17723
rect 11816 17587 11952 17723
rect 11952 17587 11956 17723
rect 11812 17583 11956 17587
rect 1614 17194 1678 17198
rect 1614 17138 1618 17194
rect 1618 17138 1674 17194
rect 1674 17138 1678 17194
rect 1614 17134 1678 17138
rect 1701 17195 1765 17199
rect 1701 17139 1705 17195
rect 1705 17139 1761 17195
rect 1761 17139 1765 17195
rect 1701 17135 1765 17139
rect 1798 17195 1942 17199
rect 1614 17114 1678 17118
rect 1614 17058 1618 17114
rect 1618 17058 1674 17114
rect 1674 17058 1678 17114
rect 1614 17054 1678 17058
rect 1701 17115 1765 17119
rect 1701 17059 1705 17115
rect 1705 17059 1761 17115
rect 1761 17059 1765 17115
rect 1701 17055 1765 17059
rect 1798 17059 1802 17195
rect 1802 17059 1938 17195
rect 1938 17059 1942 17195
rect 1798 17055 1942 17059
rect 22652 15138 22796 15142
rect 22652 15002 22656 15138
rect 22656 15002 22792 15138
rect 22792 15002 22796 15138
rect 22652 14998 22796 15002
rect 26516 14451 26660 14455
rect 26516 14315 26520 14451
rect 26520 14315 26656 14451
rect 26656 14315 26660 14451
rect 26516 14311 26660 14315
rect 232 13322 296 13326
rect 232 13266 236 13322
rect 236 13266 292 13322
rect 292 13266 296 13322
rect 232 13262 296 13266
rect 319 13323 383 13327
rect 319 13267 323 13323
rect 323 13267 379 13323
rect 379 13267 383 13323
rect 319 13263 383 13267
rect 416 13323 560 13327
rect 232 13242 296 13246
rect 232 13186 236 13242
rect 236 13186 292 13242
rect 292 13186 296 13242
rect 232 13182 296 13186
rect 319 13243 383 13247
rect 319 13187 323 13243
rect 323 13187 379 13243
rect 379 13187 383 13243
rect 319 13183 383 13187
rect 416 13187 420 13323
rect 420 13187 556 13323
rect 556 13187 560 13323
rect 416 13183 560 13187
rect 18788 13000 18932 13004
rect 18788 12864 18792 13000
rect 18792 12864 18928 13000
rect 18928 12864 18932 13000
rect 18788 12860 18932 12864
rect 22652 10784 22796 10788
rect 22652 10648 22656 10784
rect 22656 10648 22792 10784
rect 22792 10648 22796 10784
rect 22652 10644 22796 10648
rect 4948 4622 5012 4686
rect 5035 4623 5099 4687
rect 4948 4542 5012 4606
rect 5035 4543 5099 4607
rect 27569 2424 27713 2428
rect 27569 2288 27573 2424
rect 27573 2288 27709 2424
rect 27709 2288 27713 2424
rect 27569 2284 27713 2288
rect 30380 2158 30524 2162
rect 30380 2022 30384 2158
rect 30384 2022 30520 2158
rect 30520 2022 30524 2158
rect 30380 2018 30524 2022
rect 26516 1901 26660 1905
rect 26516 1765 26520 1901
rect 26520 1765 26656 1901
rect 26656 1765 26660 1901
rect 26516 1761 26660 1765
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 800 44760 26066 44952
rect 200 41540 600 44152
rect 200 41539 319 41540
rect 200 41475 232 41539
rect 296 41476 319 41539
rect 383 41476 416 41540
rect 296 41475 416 41476
rect 200 41460 416 41475
rect 200 41459 319 41460
rect 200 41395 232 41459
rect 296 41396 319 41459
rect 383 41396 416 41460
rect 560 41396 600 41540
rect 296 41395 600 41396
rect 200 22609 600 41395
rect 200 22608 319 22609
rect 200 22544 232 22608
rect 296 22545 319 22608
rect 383 22545 416 22609
rect 296 22544 416 22545
rect 200 22529 416 22544
rect 200 22528 319 22529
rect 200 22464 232 22528
rect 296 22465 319 22528
rect 383 22465 416 22529
rect 560 22465 600 22609
rect 296 22464 600 22465
rect 200 13327 600 22464
rect 200 13326 319 13327
rect 200 13262 232 13326
rect 296 13263 319 13326
rect 383 13263 416 13327
rect 296 13262 416 13263
rect 200 13247 416 13262
rect 200 13246 319 13247
rect 200 13182 232 13246
rect 296 13183 319 13246
rect 383 13183 416 13247
rect 560 13183 600 13327
rect 296 13182 600 13183
rect 200 1000 600 13182
rect 800 33793 1200 44760
rect 20734 41547 20914 41556
rect 20734 41403 20752 41547
rect 20896 41403 20914 41547
rect 20734 41392 20914 41403
rect 800 33765 2465 33793
rect 800 33764 2206 33765
rect 800 33700 2119 33764
rect 2183 33701 2206 33764
rect 2270 33701 2303 33765
rect 2183 33700 2303 33701
rect 800 33685 2303 33700
rect 800 33684 2206 33685
rect 800 33620 2119 33684
rect 2183 33621 2206 33684
rect 2270 33621 2303 33685
rect 2447 33621 2465 33765
rect 2183 33620 2465 33621
rect 800 33593 2465 33620
rect 800 17227 1200 33593
rect 11794 17727 11974 17736
rect 11794 17583 11812 17727
rect 11956 17583 11974 17727
rect 11794 17572 11974 17583
rect 800 17199 1960 17227
rect 800 17198 1701 17199
rect 800 17134 1614 17198
rect 1678 17135 1701 17198
rect 1765 17135 1798 17199
rect 1678 17134 1798 17135
rect 800 17119 1798 17134
rect 800 17118 1701 17119
rect 800 17054 1614 17118
rect 1678 17055 1701 17118
rect 1765 17055 1798 17119
rect 1942 17055 1960 17199
rect 1678 17054 1960 17055
rect 800 17027 1960 17054
rect 800 6392 1200 17027
rect 11852 15696 11912 17572
rect 20778 16033 20878 41392
rect 26558 37630 26618 45152
rect 26451 37621 26618 37630
rect 26451 37477 26464 37621
rect 26608 37477 26618 37621
rect 26451 37466 26618 37477
rect 26498 25988 26678 25997
rect 26498 25844 26516 25988
rect 26660 25844 26678 25988
rect 18770 15933 20878 16033
rect 22634 25084 22814 25093
rect 22634 24940 22652 25084
rect 22796 24940 22814 25084
rect 18770 15696 18950 15933
rect 11852 15636 18950 15696
rect 18770 13004 18950 15636
rect 18770 12860 18788 13004
rect 18932 12860 18950 13004
rect 800 6200 1532 6392
rect 800 1000 1200 6200
rect 4935 4687 5274 4711
rect 4935 4686 5035 4687
rect 4935 4622 4948 4686
rect 5012 4623 5035 4686
rect 5099 4623 5274 4687
rect 5012 4622 5274 4623
rect 4935 4607 5554 4622
rect 4935 4606 5035 4607
rect 4935 4542 4948 4606
rect 5012 4543 5035 4606
rect 5099 4562 5554 4607
rect 5099 4543 5274 4562
rect 5012 4542 5274 4543
rect 4935 4519 5274 4542
rect 5494 2273 5554 4562
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 12860
rect 22634 15142 22814 24940
rect 22634 14998 22652 15142
rect 22796 14998 22814 15142
rect 22634 10788 22814 14998
rect 22634 10644 22652 10788
rect 22796 10644 22814 10788
rect 22634 0 22814 10644
rect 26498 14455 26678 25844
rect 27110 24433 27170 45152
rect 27003 24424 27170 24433
rect 27003 24280 27016 24424
rect 27160 24280 27170 24424
rect 27003 24269 27170 24280
rect 26498 14311 26516 14455
rect 26660 14311 26678 14455
rect 26498 1905 26678 14311
rect 27662 2437 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 30362 26638 30542 26647
rect 30362 26494 30380 26638
rect 30524 26494 30542 26638
rect 30362 23701 30542 26494
rect 30362 23557 30380 23701
rect 30524 23557 30542 23701
rect 27556 2428 27723 2437
rect 27556 2284 27569 2428
rect 27713 2284 27723 2428
rect 27556 2273 27723 2284
rect 26498 1761 26516 1905
rect 26660 1761 26678 1905
rect 26498 0 26678 1761
rect 30362 2162 30542 23557
rect 30362 2018 30380 2162
rect 30524 2018 30542 2162
rect 30362 0 30542 2018
use pravindu_nilakna_sky130_opamp  pravindu_nilakna_sky130_opamp_0
timestamp 1591351771
transform 1 0 2263 0 1 26287
box -1805 0 18594 15246
use rajinthanr_opamp  rajinthanr_opamp_0
timestamp 1591351771
transform 1 0 404 0 1 25503
box 1309 -8828 18153 -2324
use lochidev_two_stage_opamp  two_stage_opamp_0
timestamp 1591351771
transform 1 0 0 0 1 0
box 1460 2381 11160 13833
<< labels >>
flabel metal4 s 22634 378 22814 658 0 FreeSans 600 0 0 0 Vp
port 53 nsew
flabel metal4 s 30362 425 30542 716 0 FreeSans 600 0 0 0 Iref
port 54 nsew
flabel metal4 s 26498 432 26678 692 0 FreeSans 600 0 0 0 Vm
port 55 nsew
flabel metal4 s 18770 423 18950 725 0 FreeSans 600 0 0 0 Vout
port 56 nsew
flabel metal4 s 200 1000 600 44152 1 FreeSans 500 0 0 0 VDPWR
port 52 nsew
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 600 90 0 0 clk
port 1 nsew
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 600 90 0 0 ena
port 2 nsew
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 600 90 0 0 rst_n
port 3 nsew
flabel metal4 s 30362 0 30542 200 0 FreeSans 1200 0 0 0 ua[0]
port 4 nsew
flabel metal4 s 26498 0 26678 200 0 FreeSans 1200 0 0 0 ua[1]
port 5 nsew
flabel metal4 s 22634 0 22814 200 0 FreeSans 1200 0 0 0 ua[2]
port 6 nsew
flabel metal4 s 18770 0 18950 200 0 FreeSans 1200 0 0 0 ua[3]
port 7 nsew
flabel metal4 s 14906 0 15086 200 0 FreeSans 1200 0 0 0 ua[4]
port 8 nsew
flabel metal4 s 11042 0 11222 200 0 FreeSans 1200 0 0 0 ua[5]
port 9 nsew
flabel metal4 s 7178 0 7358 200 0 FreeSans 1200 0 0 0 ua[6]
port 10 nsew
flabel metal4 s 3314 0 3494 200 0 FreeSans 1200 0 0 0 ua[7]
port 11 nsew
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 600 90 0 0 ui_in[0]
port 12 nsew
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 600 90 0 0 ui_in[1]
port 13 nsew
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 600 90 0 0 ui_in[2]
port 14 nsew
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 600 90 0 0 ui_in[3]
port 15 nsew
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 600 90 0 0 ui_in[4]
port 16 nsew
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 600 90 0 0 ui_in[5]
port 17 nsew
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 600 90 0 0 ui_in[6]
port 18 nsew
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 600 90 0 0 ui_in[7]
port 19 nsew
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 600 90 0 0 uio_in[0]
port 20 nsew
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 600 90 0 0 uio_in[1]
port 21 nsew
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 600 90 0 0 uio_in[2]
port 22 nsew
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 600 90 0 0 uio_in[3]
port 23 nsew
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 600 90 0 0 uio_in[4]
port 24 nsew
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 600 90 0 0 uio_in[5]
port 25 nsew
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 600 90 0 0 uio_in[6]
port 26 nsew
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 600 90 0 0 uio_in[7]
port 27 nsew
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 600 90 0 0 uio_oe[0]
port 28 nsew
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 600 90 0 0 uio_oe[1]
port 29 nsew
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 600 90 0 0 uio_oe[2]
port 30 nsew
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 600 90 0 0 uio_oe[3]
port 31 nsew
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 600 90 0 0 uio_oe[4]
port 32 nsew
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 600 90 0 0 uio_oe[5]
port 33 nsew
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 600 90 0 0 uio_oe[6]
port 34 nsew
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 600 90 0 0 uio_oe[7]
port 35 nsew
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 600 90 0 0 uio_out[0]
port 36 nsew
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 600 90 0 0 uio_out[1]
port 37 nsew
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 600 90 0 0 uio_out[2]
port 38 nsew
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 600 90 0 0 uio_out[3]
port 39 nsew
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 600 90 0 0 uio_out[4]
port 40 nsew
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 600 90 0 0 uio_out[5]
port 41 nsew
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 600 90 0 0 uio_out[6]
port 42 nsew
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 600 90 0 0 uio_out[7]
port 43 nsew
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 600 90 0 0 uo_out[0]
port 44 nsew
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 600 90 0 0 uo_out[1]
port 45 nsew
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 600 90 0 0 uo_out[2]
port 46 nsew
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 600 90 0 0 uo_out[3]
port 47 nsew
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 600 90 0 0 uo_out[4]
port 48 nsew
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 600 90 0 0 uo_out[5]
port 49 nsew
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 600 90 0 0 uo_out[6]
port 50 nsew
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 600 90 0 0 uo_out[7]
port 51 nsew
flabel metal4 s 800 1000 1200 44152 1 FreeSans 500 0 0 0 VGND
port 57 nsew
<< properties >>
string FIXED_BBOX 0 0 32180 45152
string path 93.850 79.915 104.140 79.915 104.140 207.780 
<< end >>
